// ---------------------------------------------
// Interface: coffee-if
// ---------------------------------------------
interface coffee_if(
  input logic 	clk
);
  logic 		size;
  logic			with_milk;
  logic			with_foam;
  logic [2:0]	coffee_type;
  
endinterface: coffee_if