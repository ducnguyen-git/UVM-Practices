interface our_interface(input logic clk);

	// Inputs
	logic [7:0] input_1;
	logic [7:0] input_2;
	
	// Output
	logic [15:0] output;

endinterface
